module main

import divagame

fn main() {
	divagame.run()
}
