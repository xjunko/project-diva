module enums

pub const clip_part = 1
pub const clip_all = 2

pub const command_jump = 1
pub const command_clip = 2
pub const command_rect = 3
pub const command_text = 4
pub const command_icon = 5
pub const command_max = 6

pub const color_text = 0
pub const color_border = 1
pub const color_windowbg = 2
pub const color_titlebg = 3
pub const color_titletext = 4
pub const color_panelbg = 5
pub const color_button = 6
pub const color_buttonhover = 7
pub const color_buttonfocus = 8
pub const color_base = 9
pub const color_basehover = 10
pub const color_basefocus = 11
pub const color_scrollbase = 12
pub const color_scrollthumb = 13
pub const color_max = 14
